`include "defines.sv"


module  test_utils(     input   logic       clk, reset, we,
                        input   logic [`MEM_DATA_BUS]   wd,
                        input   logic[`MEM_ADDR_BUS]    a,
                        input   logic[`MEM_WMASK_BUS]   wmask,
                        output  logic[`MEM_DATA_BUS]    rd);
        logic [`MEM_DATA_BUS]   begin_signature
endmodule
