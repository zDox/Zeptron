module datapath();
endmodule
