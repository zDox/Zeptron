`include "defines.sv"

module execution_stage(// Inputs from General
                        input   logic                   clk, reset,
                        // Inputs from ID
                        input   logic [`INSTR_BUS]      instr, pc,
                        controlsgs_if                   controls,
                        // Inputs from WB
                        input   logic                   regwe,
                        input   logic [`REG_ADDR_BUS]   regwa,
                        input   logic [`REG_BUS]        regwd,
                        // Output to IF and DM
                        output  logic [`MEM_DATA_BUS]   alu_y,
                        // Outputs to DM
                        output  logic [`MEM_DATA_BUS]   rdd2,
                        output  logic [`REG_ADDR_BUS]   rd,
                        // Outputs to IF
                        output  logic [`INSTR_ADDR_BUS] pc_4,
                        output  logic                   b_taken);
    logic [`REG_ADDR_BUS]   rs1, rs2;
    logic [`REG_BUS]        rrd1, imm;
    logic [`REG_BUS]        srca, srcb;

    // Determine rs1 and rs2
    assign rs1 = instr[19:15];
    assign rs2 = instr[24:20];

    register_file       reg_file(   .clk(clk), .reset(reset),
                                    .ra1(rs1), .ra2(rs2),
                                    .wa3(regwa), .wd3(regwd), .we3(regwe),
                                    .rd1(rrd1), .rd2(rrd2));
    immediate_generator ig (        .instr(instr), .y(imm));


    // ALU
    mux4                mux_srca(   .d1(rrd1), .d2({32{1'b0}}), .d3(pc), .y(srca));
    mux2                mux_srcb(   .d1(rrd2), .d2(imm), .y(srcb));
    alu                 alu(        .a(srca), .b(srcb), .alu_op(controls.alu_op),
                                    .y(alu_y));

    jump_control        jc(         .bj_op(controls.bj_op),
                                    .srca(srca), .srcb(srcb),
                                    .b_taken(b_taken));

    // PC_4 and PC_IMM calculation
    adder               add_pc4(    .a(pc), .b(4), .y(pc_4));
endmodule
