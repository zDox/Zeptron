module alu(input    logic [31:0]    a, b,
           input    logic [3:0]     aluop,
           output   logic [31:0]    y,
           output   logic           z);

endmodule
