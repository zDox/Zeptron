module riscv ();
endmodule
