module controller();
endmodule
