module sign_extension(  input   logic [31:0] a,
                        output  logic [31:0] y);
endmodule
